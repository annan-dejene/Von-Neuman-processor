// `include "ALU.v"
// `include "regfile.v"
// `include "pc.v"
// `include "control_unit.v"

module datapath(clock, reset, instruction_register, pc_write_enable, mem_read_data_in, instruction_address, mem_write_enable_out, mem_address_select_out, mem_write_data_out, alu_address_out, halt_cpu_out);
    input clock;
    input reset;
    input [15:0] instruction_register; // Instruction coming from memory
    output [7:0] instruction_address;  // PC address to memory module

    input wire [15:0] mem_read_data_in;

    // NEW: Input to freeze the PC when needed
    input pc_write_enable; 
    
 
    // NEW PORTS ADDED FOR TOP-LEVEL MEMORY CONTROL:
    output wire mem_write_enable_out;
    output wire mem_address_select_out;
    output wire [15:0] mem_write_data_out; // Data to write to memory
    output wire [7:0] alu_address_out;      // Address to write/read from memory (ALU result)
    output wire halt_cpu_out;   // Halt signal to stop simulation


    // --------------------------------------------------
    // Internal Wires for the Control Signals (Generated by Control Unit, defined here)
    // We instantiate them as wires here, the control unit module will drive them later.
    // --------------------------------------------------
    wire reg_write_enable_ctrl;
    wire mem_write_enable_ctrl;
    wire [3:0] alu_opcode_ctrl; 
    wire alu_src_select_ctrl;       // 0: Use RegFile data2, 1: Use Immediate value depending on the instruction type ----> set by the control unit
    wire mem_to_reg_select_ctrl;    // 0: Write ALU result to RegFile, 1: Write Memory data to RegFile
    // Add other control signals as needed (e.g., jump enable, halt enable)
    wire halt_cpu_ctrl;
    wire jump_enable_ctrl;
    wire branch_enable_ctrl; // declared here so it's visible and can be connected to the top-level outputs

    wire mem_address_select_ctrl;

    // --------------------------------------------------
    // Internal Wires for Data Flow
    // --------------------------------------------------
    wire [7:0] pc_next_address; // PC address calculated (PC+1, branch target, or jump target)
    wire [15:0] regfile_data1_out, regfile_data2_out; // Outputs from RegFile --> content of the selected registers
    wire [15:0] alu_result_out;
    wire alu_zero_flag;

    // --------------------------------------------------
    // Instruction Decoding Wires (based on your ISA format) --- decoded from the instruction register
    // --------------------------------------------------
    wire [3:0] opcode;
    wire [2:0] rd_addr, rs_addr, rt_addr;
    wire [5:0] immediate;

    assign opcode = instruction_register[15:12];
    assign rd_addr = instruction_register[11:9];
    assign rs_addr = instruction_register[8:6];
    assign rt_addr = instruction_register[5:3];
    assign immediate = instruction_register[5:0]; // The immediate is 6 bits for I-type format instructions --------

// ----> we wil use either rs and rt for R-type instructions or the immediate 9 bits for I-type instructions
    
    // We need to sign-extend the 6-bit immediate to 16 bits for arithmetic operations (MOV, LD, ST, BEQZ)
    wire [15:0] immediate_sign_extended;
    assign immediate_sign_extended = {{10{immediate[5]}}, immediate}; // Sign extend 6 bits to 16 bits

    // --------------------------------------------------
    // MUXes and Logic
    // --------------------------------------------------

    // MUX 1: ALU Source B selection (RegFile data2 or immediate value)
    wire [15:0] regfile_immediate_mux_ALU;

    assign regfile_immediate_mux_ALU = (alu_src_select_ctrl == 0) ? regfile_data2_out : immediate_sign_extended;


    // MUX 2: Register File Write Data Selection (ALU result or Memory Read Data)
    wire [15:0] reg_write_data_in;
    assign reg_write_data_in = (mem_to_reg_select_ctrl == 0) ? alu_result_out : mem_read_data_in;


    // --------------------------------------------------
    // PC Control Logic & MUXes (for sequential, branch, jump) - FIX 1 APPLIED
    // --------------------------------------------------
    wire [7:0] pc_plus_1;
    assign pc_plus_1 = instruction_address + 8'd1;

    // Calculate Branch Target Address: PC+1 + offset (sign extended)
    // Note: The result needs to be trimmed to 8 bits for your 8-bit address space
    wire [7:0] branch_target_address;
    assign branch_target_address = immediate_sign_extended[7:0]; 
    
    // For JMP (OP_JMP), we use the immediate value as the target address (absolute address)
    wire [7:0] pc_jump_target;
    assign pc_jump_target = immediate_sign_extended[7:0]; 

    // MUX 3 (PC Source MUX): 
    // Uses priority encoding: Jump > Branch Taken > PC+1
    assign pc_next_address = (jump_enable_ctrl) ? pc_jump_target : 
                                                                    (branch_enable_ctrl && alu_zero_flag) ? branch_target_address : pc_plus_1;                                 

    // --------------------------------------------------
    // PC Logic with Stall (Write Enable)
    // --------------------------------------------------
    // If pc_write_enable is 0, we force the "next" address to be the "current" address.
    // This effectively holds the PC value for one cycle.
    // We need to do this to be able to fetch data or store data to memory while the program counter is frozen and not incremented as we are unable to fetch next instruction and data from the same memory with the same data path i.e. the von neumann bottle neck
    wire [7:0] actual_next_pc;
    assign actual_next_pc = (pc_write_enable) ? pc_next_address : instruction_address;



    // --------------------------------------------------
    // Component Instantiations (PC, Regfile, ALU)
    // --------------------------------------------------

    // Program Counter (pc)
    pc my_pc(
        .clock(clock),
        .reset(reset),
        .next_address(actual_next_pc), // Simple sequential increment for now
        .current_address(instruction_address)
    );

    // Register File (regfile)
    regfile my_regfile(
        .regSource1(rs_addr),
        .regSource2(rt_addr),
        .regDestination(rd_addr), // Destination address comes from the instruction [11:9]
        .writeData(reg_write_data_in),
        .data1(regfile_data1_out),
        .data2(regfile_data2_out),
        .writeEnable(reg_write_enable_ctrl && pc_write_enable),
        .clock(clock),
        .reset(reset)
    );

    // Instantiate ALU (ALU)
    ALU my_alu(
        .num1(regfile_data1_out),
        .num2(regfile_immediate_mux_ALU),
        .opcode(alu_opcode_ctrl),
        .result(alu_result_out),
        .zero(alu_zero_flag)
    );

    // --------------------------------------------------
    // Connect internal control/data wires to module outputs so top-level can use them
    // --------------------------------------------------
    // Drive memory control/data outputs
    // During reset ensure safe defaults so memory fetch can use PC (no dependence on decoded opcode)
    assign mem_write_enable_out = reset ? 1'b0 : mem_write_enable_ctrl;
    assign mem_address_select_out = reset ? 1'b0 : mem_address_select_ctrl;
    assign mem_write_data_out = reset ? 16'h0000 : regfile_data2_out; // write data comes from regfile data2
    assign alu_address_out = reset ? 8'h00 : alu_result_out[7:0];   // lower 8 bits of ALU result used as memory address
    assign halt_cpu_out = reset ? 1'b0 : halt_cpu_ctrl;
    

    // --------------------------------------------------
    // Control Unit Instantiation
    // --------------------------------------------------
    // Connect the control unit to all our new wires/signals
    control_unit my_control_unit(
        .opcode(opcode),
        .alu_zero_flag_in(alu_zero_flag),
        .reg_write_enable_out(reg_write_enable_ctrl), // write enabe for register file ---> set to 1 when writing to register file
        .mem_write_enable_out(mem_write_enable_ctrl), // write enable for memory ----> set to 1 when writing to memory
        .alu_opcode_out(alu_opcode_ctrl), // the opcode for the ALU operation outputted from the control unit based on the instruction register[15:12] and inputted to the ALU instance to select operation
        .alu_src_select_out(alu_src_select_ctrl), //set by the control unit as output depending on the instruction whether it uses register file data 2 or immediate --> 0: Use RegFile data2, 1: Use Immediate value depending on the instruction type 
        .mem_to_reg_select_out(mem_to_reg_select_ctrl), // 0: Write ALU result to RegFile, 1: Write Memory data to RegFile
        .halt_cpu_out(halt_cpu_ctrl),
        .jump_enable_out(jump_enable_ctrl),
        .branch_enable_out(branch_enable_ctrl), // Connect new control signal
        .mem_address_select_out(mem_address_select_ctrl) // Connect new control signal
    );


endmodule
