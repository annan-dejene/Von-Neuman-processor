`include "ALU.v"
`include "regfile.v"
`include "pc.v"
`include "control_unit.v"

module datapath(clock, reset, instruction_address, instruction_register, mem_write_enable_out, mem_address_select_out, mem_write_data_out, alu_address_out, halt_cpu_out);
    input clock;
    input reset;
    output [7:0] instruction_address;  // PC address to memory module
    input [15:0] instruction_register; // Instruction coming from memory

    // NEW PORTS ADDED FOR TOP-LEVEL MEMORY CONTROL:
    output wire mem_write_enable_out;
    output wire mem_address_select_out;
    output wire [15:0] mem_write_data_out; // Data to write to memory
    output wire [7:0] alu_address_out;      // Address to write/read from memory (ALU result)
    output wire halt_cpu_out;   // Halt signal to stop simulation


    // --------------------------------------------------
    // Internal Wires for the Control Signals (Generated by Control Unit, defined here)
    // We instantiate them as wires here, the control unit module will drive them later.
    // --------------------------------------------------
    wire reg_write_enable_ctrl;
    wire mem_write_enable_ctrl;
    wire [3:0] alu_opcode_ctrl; 
    wire alu_src_select_ctrl;       // 0: Use RegFile data2, 1: Use Immediate value depending on the instruction type ----> set by the control unit
    wire mem_to_reg_select_ctrl;    // 0: Write ALU result to RegFile, 1: Write Memory data to RegFile
    // Add other control signals as needed (e.g., jump enable, halt enable)
    wire halt_cpu_ctrl;
    wire jump_enable_ctrl;


    // --------------------------------------------------
    // Internal Wires for Data Flow
    // --------------------------------------------------
    wire [7:0] pc_next_address; // PC address calculated (PC+1, branch target, or jump target)
    wire [15:0] regfile_data1_out, regfile_data2_out; // Outputs from RegFile --> content of the selected registers
    wire [15:0] alu_result_out;
    wire alu_zero_flag;

    // --------------------------------------------------
    // Instruction Decoding Wires (based on your ISA format) --- decoded from the instruction register
    // --------------------------------------------------
    wire [3:0] opcode;
    wire [2:0] rd_addr, rs_addr, rt_addr;
    wire [5:0] immediate;

    assign opcode = instruction_register[15:12];
    assign rd_addr = instruction_register[11:9];
    assign rs_addr = instruction_register[8:6];
    assign rt_addr = instruction_register[5:3];
    assign immediate = instruction_register[5:0]; // The immediate is 6 bits for I-type format instructions --------

// ----> we wil use either rs and rt for R-type instructions or the immediate 9 bits for I-type instructions
    
    // We need to sign-extend the 6-bit immediate to 16 bits for arithmetic operations (MOV, LD, ST, BEQZ)
    wire [15:0] immediate_sign_extended;
    assign immediate_sign_extended = {{10{immediate[5]}}, immediate}; // Sign extend 6 bits to 16 bits

    // --------------------------------------------------
    // MUXes and Logic
    // --------------------------------------------------

    // MUX 1: ALU Source B selection (RegFile data2 or immediate value)
    wire [15:0] regfile_immediate_mux_ALU;

    assign regfile_immediate_mux_ALU = (alu_src_select_ctrl == 0) ? regfile_data2_out : immediate_sign_extended;


    // MUX 2: Register File Write Data Selection (ALU result or Memory Read Data)
    wire [15:0] reg_write_data_in;
    assign reg_write_data_in = (mem_to_reg_select_ctrl == 0) ? alu_result_out : mem_read_data_out;


    // --------------------------------------------------
    // PC Control Logic & MUXes (for sequential, branch, jump) - FIX 1 APPLIED
    // --------------------------------------------------
    wire [7:0] pc_plus_1;
    assign pc_plus_1 = instruction_address + 8'd1;

    // Calculate Branch Target Address: PC+1 + offset (sign extended)
    // Note: The result needs to be trimmed to 8 bits for your 8-bit address space
    wire [7:0] branch_target_address;
    assign branch_target_address = instruction_address + immediate_sign_extended[7:0] + 8'd1; 
    
    // For JMP (OP_JMP), we use the immediate value as the target address (absolute address)
    wire [7:0] pc_jump_target;
    assign pc_jump_target = immediate_sign_extended[7:0]; 

    // MUX 3 (PC Source MUX): 
    // Uses priority encoding: Jump > Branch Taken > PC+1
    assign pc_next_address = (jump_enable_ctrl) ? pc_jump_target : 
                                                                    (branch_enable_ctrl && alu_zero_flag) ? branch_target_address : pc_plus_1;                                 


    // --------------------------------------------------
    // Component Instantiations (PC, Regfile, ALU)
    // --------------------------------------------------

    // Program Counter (pc)
    pc my_pc(
        .clock(clock),
        .reset(reset),
        .next_address(pc_next_address), // Simple sequential increment for now
        .current_address(instruction_address)
    );

    // Register File (regfile)
    regfile my_regfile(
        .regSource1(rs_addr),
        .regSource2(rt_addr),
        .regDestination(rd_addr), // Destination address comes from the instruction [11:9]
        .writeData(reg_write_data_in),
        .data1(regfile_data1_out),
        .data2(regfile_data2_out),
        .writeEnable(reg_write_enable_ctrl),
        .clock(clock),
        .reset(reset)
    );

    // Instantiate ALU (ALU)
    ALU my_alu(
        .num1(regfile_data1_out),
        .num2(regfile_immediate_mux_ALU),
        .opcode(alu_opcode_ctrl),
        .result(alu_result_out),
        .zero(alu_zero_flag)
    );
    

    // --------------------------------------------------
    // Control Unit Instantiation
    // --------------------------------------------------
    // Connect the control unit to all our new wires/signals
    control_unit my_control_unit(
        .opcode(opcode),
        .alu_zero_flag_in(alu_zero_flag),
        .reg_write_enable_out(reg_write_enable_ctrl),
        .mem_write_enable_out(mem_write_enable_ctrl),
        .alu_opcode_out(alu_opcode_ctrl),
        .alu_src_select_out(alu_src_select_ctrl),
        .mem_to_reg_select_out(mem_to_reg_select_ctrl),
        .halt_cpu_out(halt_cpu_ctrl),
        .jump_enable_out(jump_enable_ctrl),
        .branch_enable_out(branch_enable_ctrl), // Connect new control signal
        .mem_address_select_out(mem_address_select_ctrl) // Connect new control signal
    );


endmodule
